/*
    pe集群控制模块。我们需要将其用有限状态机进行控制，复用pe集群。
    状态1:  IDLE。该状态下所有的寄存器的值都应该归零。从磁盘中读入数据，存储在寄存器中准备进行运算。
    状态2:  SELF。自注意力第一步。我们需要将8x4的矩阵和4x8的矩阵相乘得到8x8的矩阵，并进行量化后存储。
            随后在每一列（行）完成运算后
*/
`include "pe_8x8_cluster.v"
module pe_8x8_top(

);
endmodule